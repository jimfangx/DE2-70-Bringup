library verilog;
use verilog.vl_types.all;
entity tb_reset_delay is
end tb_reset_delay;
