library verilog;
use verilog.vl_types.all;
entity tb_BasicTests is
end tb_BasicTests;
