library verilog;
use verilog.vl_types.all;
entity tb_VGA_Controller is
end tb_VGA_Controller;
