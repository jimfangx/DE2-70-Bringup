library verilog;
use verilog.vl_types.all;
entity tb_VGA is
end tb_VGA;
